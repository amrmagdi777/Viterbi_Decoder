library verilog;
use verilog.vl_types.all;
entity branch_metric is
    generic(
        S1              : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        S2              : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        S3              : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        S4              : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi1);
        S5              : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        S6              : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi1);
        S7              : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        S8              : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        state1_1_output : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        state1_2_output : vl_logic_vector(0 to 1) := (Hi1, Hi1);
        state2_4_output : vl_logic_vector(0 to 1) := (Hi0, Hi1);
        state2_3_output : vl_logic_vector(0 to 1) := (Hi1, Hi0);
        state3_5_output : vl_logic_vector(0 to 1) := (Hi0, Hi1);
        state3_6_output : vl_logic_vector(0 to 1) := (Hi1, Hi0);
        state4_8_output : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        state4_7_output : vl_logic_vector(0 to 1) := (Hi1, Hi1);
        state5_2_output : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        state5_1_output : vl_logic_vector(0 to 1) := (Hi1, Hi1);
        state6_3_output : vl_logic_vector(0 to 1) := (Hi0, Hi1);
        state6_4_output : vl_logic_vector(0 to 1) := (Hi1, Hi0);
        state7_5_output : vl_logic_vector(0 to 1) := (Hi1, Hi0);
        state7_6_output : vl_logic_vector(0 to 1) := (Hi0, Hi1);
        state8_7_output : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        state8_8_output : vl_logic_vector(0 to 1) := (Hi1, Hi1)
    );
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        sys             : in     vl_logic;
        parity          : in     vl_logic;
        branch_enable   : in     vl_logic;
        state1_1_error  : out    vl_logic_vector(1 downto 0);
        state1_2_error  : out    vl_logic_vector(1 downto 0);
        state2_4_error  : out    vl_logic_vector(1 downto 0);
        state2_3_error  : out    vl_logic_vector(1 downto 0);
        state3_5_error  : out    vl_logic_vector(1 downto 0);
        state3_6_error  : out    vl_logic_vector(1 downto 0);
        state4_8_error  : out    vl_logic_vector(1 downto 0);
        state4_7_error  : out    vl_logic_vector(1 downto 0);
        state5_2_error  : out    vl_logic_vector(1 downto 0);
        state5_1_error  : out    vl_logic_vector(1 downto 0);
        state6_3_error  : out    vl_logic_vector(1 downto 0);
        state6_4_error  : out    vl_logic_vector(1 downto 0);
        state7_6_error  : out    vl_logic_vector(1 downto 0);
        state7_5_error  : out    vl_logic_vector(1 downto 0);
        state8_7_error  : out    vl_logic_vector(1 downto 0);
        state8_8_error  : out    vl_logic_vector(1 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of S1 : constant is 1;
    attribute mti_svvh_generic_type of S2 : constant is 1;
    attribute mti_svvh_generic_type of S3 : constant is 1;
    attribute mti_svvh_generic_type of S4 : constant is 1;
    attribute mti_svvh_generic_type of S5 : constant is 1;
    attribute mti_svvh_generic_type of S6 : constant is 1;
    attribute mti_svvh_generic_type of S7 : constant is 1;
    attribute mti_svvh_generic_type of S8 : constant is 1;
    attribute mti_svvh_generic_type of state1_1_output : constant is 1;
    attribute mti_svvh_generic_type of state1_2_output : constant is 1;
    attribute mti_svvh_generic_type of state2_4_output : constant is 1;
    attribute mti_svvh_generic_type of state2_3_output : constant is 1;
    attribute mti_svvh_generic_type of state3_5_output : constant is 1;
    attribute mti_svvh_generic_type of state3_6_output : constant is 1;
    attribute mti_svvh_generic_type of state4_8_output : constant is 1;
    attribute mti_svvh_generic_type of state4_7_output : constant is 1;
    attribute mti_svvh_generic_type of state5_2_output : constant is 1;
    attribute mti_svvh_generic_type of state5_1_output : constant is 1;
    attribute mti_svvh_generic_type of state6_3_output : constant is 1;
    attribute mti_svvh_generic_type of state6_4_output : constant is 1;
    attribute mti_svvh_generic_type of state7_5_output : constant is 1;
    attribute mti_svvh_generic_type of state7_6_output : constant is 1;
    attribute mti_svvh_generic_type of state8_7_output : constant is 1;
    attribute mti_svvh_generic_type of state8_8_output : constant is 1;
end branch_metric;
